/**
 * Author: Borys Strzebonski
 *
 * Description:
 * Bitmaps for letters (simple 5x7 font)
 */

logic [6:0][4:0] letter_E = '{
    5'b11111,
    5'b00001,
    5'b00001,
    5'b11111,
    5'b00001,
    5'b00001,
    5'b11111
};

logic [6:0][4:0] letter_A = '{
    5'b01110,
    5'b10001,
    5'b10001,
    5'b11111,
    5'b10001,
    5'b10001,
    5'b10001
};

logic [6:0][4:0] letter_L = '{
    5'b00001,
    5'b00001,
    5'b00001,
    5'b00001,
    5'b00001,
    5'b00001,
    5'b11111
};

logic [6:0][4:0] letter_H = '{
    5'b10001,
    5'b10001,
    5'b10001,
    5'b11111,
    5'b10001,
    5'b10001,
    5'b10001
};

logic [6:0][4:0] letter_I = '{
    5'b11111,
    5'b00100,
    5'b00100,
    5'b00100,
    5'b00100,
    5'b00100,
    5'b11111
};

logic [6:0][4:0] letter_T = '{
    5'b11111,
    5'b00100,
    5'b00100,
    5'b00100,
    5'b00100,
    5'b00100,
    5'b00100
};

logic [6:0][4:0] letter_S = '{
    5'b11110,
    5'b00001,
    5'b00001,
    5'b11110,
    5'b10000,
    5'b10000,
    5'b01111
};

logic [6:0][4:0] letter_N = '{
    5'b10001,
    5'b10011,
    5'b10101,
    5'b11001,
    5'b10001,
    5'b10001,
    5'b10001
};

logic [6:0][4:0] letter_D = '{
    5'b01111,
    5'b10001,
    5'b10001,
    5'b10001,
    5'b10001,
    5'b10001,
    5'b01111
};

