module char_16x16(
        input wire clk,
        input logic [7:0] char_xy,
        output logic [6:0] char_code
    );
    logic [6:0] data;

    always_ff @(posedge clk)
        char_code <= data;

    always_comb begin
        case(char_xy)
            8'h00: data = "L";
            8'h01: data = "I";
            8'h02: data = "T";
            8'h03: data = "W";
            8'h04: data = "O";
            8'h05: data = " ";
            8'h06: data = "O";
            8'h07: data = "J";
            8'h08: data = "C";
            8'h09: data = "Z";
            8'h0a: data = "Y";
            8'h0b: data = "Z";
            8'h0c: data = "N";
            8'h0d: data = "O";
            8'h0e: data = " ";
            8'h0f: data = "M";
            8'h10: data = "O";
            8'h11: data = "J";
            8'h12: data = "A";
            8'h13: data = " ";
            8'h14: data = "T";
            8'h15: data = "Y";
            8'h16: data = " ";
            8'h17: data = "J";
            8'h18: data = "E";
            8'h19: data = "S";
            8'h1a: data = "T";
            8'h1b: data = "E";
            8'h1c: data = "S";
            8'h1d: data = " ";
            8'h1e: data = "J";
            8'h1f: data = "A";
            8'h20: data = "K";
            8'h21: data = " ";
            8'h22: data = "Z";
            8'h23: data = "D";
            8'h24: data = "R";
            8'h25: data = "O";
            8'h26: data = "W";
            8'h27: data = "I";
            8'h28: data = "E";
            8'h29: data = " ";
            8'h2a: data = "I";
            8'h2b: data = "L";
            8'h2c: data = "E";
            8'h2d: data = " ";
            8'h2e: data = "C";
            8'h2f: data = "I";
            8'h30: data = "E";
            8'h31: data = " ";
            8'h32: data = "T";
            8'h33: data = "R";
            8'h34: data = "Z";
            8'h35: data = "E";
            8'h36: data = "B";
            8'h37: data = "A";
            8'h38: data = " ";
            8'h39: data = "C";
            8'h3a: data = "E";
            8'h3b: data = "N";
            8'h3c: data = "I";
            8'h3d: data = "C";
            8'h3e: data = " ";
            8'h3f: data = "T";
            8'h40: data = "E";
            8'h41: data = "N";
            8'h42: data = " ";
            8'h43: data = "T";
            8'h44: data = "Y";
            8'h45: data = "L";
            8'h46: data = "K";
            8'h47: data = "O";
            8'h48: data = " ";
            8'h49: data = "S";
            8'h4a: data = "I";
            8'h4b: data = "E";
            8'h4c: data = " ";
            8'h4d: data = "D";
            8'h4e: data = "O";
            8'h4f: data = "W";
            8'h50: data = "I";
            8'h51: data = "E";
            8'h52: data = " ";
            8'h53: data = "K";
            8'h54: data = "T";
            8'h55: data = "O";
            8'h56: data = " ";
            8'h57: data = "C";
            8'h58: data = "I";
            8'h59: data = "E";
            8'h5a: data = " ";
            8'h5b: data = "S";
            8'h5c: data = "T";
            8'h5d: data = "R";
            8'h5e: data = "A";
            8'h5f: data = "C";
            8'h60: data = "I";
            8'h61: data = "L";
            8'h62: data = " ";
            8'h63: data = "D";
            8'h64: data = "Z";
            8'h65: data = "I";
            8'h66: data = "S";
            8'h67: data = " ";
            8'h68: data = "P";
            8'h69: data = "I";
            8'h6a: data = "E";
            8'h6b: data = "K";
            8'h6c: data = "N";
            8'h6d: data = "O";
            8'h6e: data = "S";
            8'h6f: data = "C";
            8'h70: data = " ";
            8'h71: data = "T";
            8'h72: data = "W";
            8'h73: data = "A";
            8'h74: data = " ";
            8'h75: data = "W";
            8'h76: data = " ";
            8'h77: data = "C";
            8'h78: data = "A";
            8'h79: data = "L";
            8'h7a: data = "E";
            8'h7b: data = "J";
            8'h7c: data = " ";
            8'h7d: data = "O";
            8'h7e: data = "Z";
            8'h7f: data = "D";
            8'h80: data = "O";
            8'h81: data = "B";
            8'h82: data = "I";
            8'h83: data = "E";
            8'h84: data = " ";
            8'h85: data = "W";
            8'h86: data = "I";
            8'h87: data = "D";
            8'h88: data = "Z";
            8'h89: data = "E";
            8'h8a: data = " ";
            8'h8b: data = "I";
            8'h8c: data = " ";
            8'h8d: data = "O";
            8'h8e: data = "P";
            8'h8f: data = "I";
            8'h90: data = "S";
            8'h91: data = "U";
            8'h92: data = "J";
            8'h93: data = "E";
            8'h94: data = " ";
            8'h95: data = "B";
            8'h96: data = "O";
            8'h97: data = " ";
            8'h98: data = "T";
            8'h99: data = "E";
            8'h9a: data = "S";
            8'h9b: data = "K";
            8'h9c: data = "N";
            8'h9d: data = "I";
            8'h9e: data = "E";
            8'h9f: data = " ";
            8'ha0: data = "P";
            8'ha1: data = "O";
            8'ha2: data = " ";
            8'ha3: data = "T";
            8'ha4: data = "O";
            8'ha5: data = "B";
            8'ha6: data = "I";
            8'ha7: data = "E";
            8'ha8: data = " ";
            8'ha9: data = " ";
            8'haa: data = " ";
            8'hab: data = " ";
            8'hac: data = " ";
            8'had: data = " ";
            8'hae: data = " ";
            8'haf: data = " ";
            8'hb0: data = " ";
            8'hb1: data = "N";
            8'hb2: data = "A";
            8'hb3: data = "M";
            8'hb4: data = " ";
            8'hb5: data = "S";
            8'hb6: data = "T";
            8'hb7: data = "R";
            8'hb8: data = "Z";
            8'hb9: data = "E";
            8'hba: data = "L";
            8'hbb: data = "A";
            8'hbc: data = "C";
            8'hbd: data = " ";
            8'hbe: data = "N";
            8'hbf: data = "I";
            8'hc0: data = "E";
            8'hc1: data = " ";
            8'hc2: data = "K";
            8'hc3: data = "A";
            8'hc4: data = "Z";
            8'hc5: data = "A";
            8'hc6: data = "N";
            8'hc7: data = "O";
            8'hc8: data = " ";
            8'hc9: data = "W";
            8'hca: data = "S";
            8'hcb: data = "T";
            8'hcc: data = "A";
            8'hcd: data = "P";
            8'hce: data = "I";
            8'hcf: data = "L";
            8'hd0: data = "E";
            8'hd1: data = "M";
            8'hd2: data = " ";
            8'hd3: data = "N";
            8'hd4: data = "A";
            8'hd5: data = " ";
            8'hd6: data = "D";
            8'hd7: data = "Z";
            8'hd8: data = "I";
            8'hd9: data = "A";
            8'hda: data = "L";
            8'hdb: data = "O";
            8'hdc: data = " ";
            8'hdd: data = "I";
            8'hde: data = " ";
            8'hdf: data = "S";
            8'he0: data = "P";
            8'he1: data = "O";
            8'he2: data = "J";
            8'he3: data = "R";
            8'he4: data = "Z";
            8'he5: data = "A";
            8'he6: data = "L";
            8'he7: data = "E";
            8'he8: data = "M";
            8'he9: data = " ";
            8'hea: data = "N";
            8'heb: data = "A";
            8'hec: data = " ";
            8'hed: data = "P";
            8'hee: data = "O";
            8'hef: data = "L";
            8'hf0: data = "E";
            8'hf1: data = " ";
            8'hf2: data = "D";
            8'hf3: data = "W";
            8'hf4: data = "I";
            8'hf5: data = "E";
            8'hf6: data = "S";
            8'hf7: data = "C";
            8'hf8: data = "I";
            8'hf9: data = "E";
            8'hfa: data = " ";
            8'hfb: data = "A";
            8'hfc: data = "R";
            8'hfd: data = "M";
            8'hfe: data = "A";
            8'hff: data = "T";
        endcase
    end
endmodule